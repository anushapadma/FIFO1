class fifo_sequence extends uvm_sequence#(fifo_seq_item);
  `uvm_object_utils(fifo_sequence)
  
  function new(string name = "fifo_sequence");
    super.new(name);
  endfunction
  
  virtual task body();
    `uvm_info(get_type_name(), $sformatf("******** Generate 16 Write REQs ********"), UVM_LOW)
    repeat(10) begin
      req =  fifo_seq_item::type_id::create("req");
      start_item(req);
      assert(req.randomize() with {i_wren == 1;});
      finish_item(req);
    end
    #10
    `uvm_info(get_type_name(), $sformatf("******** Generate 16 Read REQs ********"), UVM_LOW)
    repeat(10) begin
      req =  fifo_seq_item::type_id::create("req");
      start_item(req);
      assert(req.randomize() with { i_rden == 1;});
      finish_item(req);
    end
    #10
    `uvm_info(get_type_name(), $sformatf("******** Generate 20 Random REQs ********"), UVM_LOW)
    repeat(20) begin
      req =  fifo_seq_item::type_id::create("req");
      start_item(req);
      assert(req.randomize());
      finish_item(req);
    end
  endtask
  
endclass
  
  
